@00080000
27 05 19 56 CE E7 E6 B3 56 89 4B 8F 00 00 00 18 
00 08 00 00 00 00 01 00 68 3B 1D B6 05 15 01 00 
73 70 69 5F 69 6D 61 67 65 2E 75 62 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
18 00 00 00 18 60 DE AD A8 63 BE EF 15 00 00 02 
15 00 00 01 15 00 00 00 
