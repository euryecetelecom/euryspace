-------------------------------
---- Project: EurySPACE CCSDS RX/TX with wishbone interface
---- Design Name: ccsds_rxtx_constants
---- Version: 1.0.0
---- Description:
---- TO BE DONE
-------------------------------
---- Author(s):
---- Guillaume Rembert
-------------------------------
---- Licence:
---- MIT
-------------------------------

package ccsds_rxtx_constants is
	constant RXTX_CST: integer := 1; -- DUMMY USELESS CONSTANT
end ccsds_rxtx_constants;
